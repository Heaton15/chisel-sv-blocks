//https://www.youtube.com/watch?v=9yo3yhUijQs

/*
*
  * 1. Register File (stores RISCV Registers). If not valid, stores ROB entry id
  * 2. If ROB entry ID is found, go to ROB and grab the information that is missing
  * 3. We also could forward the results if it is immediately available
*/
module reorder_buffer #() ();
endmodule
