module prio_arbiter_lsb_to_msb(/*AUTOARG*/);
endmodule
