module sync_fifo(/*AUTOARG*/);


endmodule


module tb;
endmodule
