module skid_buffer (/*AUTOARG*/);

endmodule

module tb;
endmodule
