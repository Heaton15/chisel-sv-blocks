module async_fifo(/*AUTOARG*/);


endmodule


module tb;
endmodule
