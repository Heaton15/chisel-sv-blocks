//https://www.youtube.com/watch?v=9yo3yhUijQs
