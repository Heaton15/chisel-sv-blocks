task automatic dump(string file);
  $dumpfile(file);
  $dumpvars(0, "tb");
endtask
