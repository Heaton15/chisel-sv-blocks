module circular_buffer(/*AUTOARG*/);
endmodule

module tb;
endmodule
